// Operand bit-width
`ifndef OWIDTH
	`define OWIDTH 8'd8
`endif

// Accumulator bit-width
`ifndef AWIDTH
	`define AWIDTH 8'd27
`endif